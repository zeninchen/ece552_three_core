module branch_decoder (
    input  wire [2:0] funct3,
    input  wire is_branch,
    input wire eq,
    input wire slt,
    output wire        b_sel
);
    //TODO
endmodule