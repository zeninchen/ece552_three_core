module branch_decoder (
    input  wire [2:0] funct3,
    input  wire is_branch,
    output wire        b_sel
);

endmodule